module main

const (
	executable_path = "app.exe"
	uninstaller = $embed_file("uninstaller.exe")
)
