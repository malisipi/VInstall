module vinstall

fn C.ShellExecute(int, &u16, &u16, &u16, &u16, int)
