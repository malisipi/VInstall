module vinstall

#include <unistd.h>
fn C.geteuid() int
