module main

const (
	executable_path = "app.out"
	uninstaller = $embed_file("uninstaller.out")
)
