module main

import malisipi.vinstall

fn main(){
	vinstall.uninstall()
}
